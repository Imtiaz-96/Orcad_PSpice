* C:\Users\ASADULLAH\Documents\scamatic3-4.sch

* Schematics Version 9.2
* Sat Nov 04 12:18:10 2017



** Analysis setup **
.tran 100ns 50us
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "scamatic3-4.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
