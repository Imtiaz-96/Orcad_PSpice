* C:\Users\ASADULLAH\Documents\Schematicelectronics2.sch

* Schematics Version 9.2
* Sat Sep 16 02:25:52 2017



** Analysis setup **
.tran 0ns 5m 0 1u
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Schematicelectronics2.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
