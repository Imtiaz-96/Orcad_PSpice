* C:\Users\ASADULLAH\Documents\222fig3.sch

* Schematics Version 9.2
* Sun Jan 21 23:01:15 2018



** Analysis setup **
.TEMP 50
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "222fig3.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
