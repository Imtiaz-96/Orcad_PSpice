* C:\Users\ASADULLAH\Documents\cc112.sch

* Schematics Version 9.2
* Tue Aug 29 08:30:47 2017



** Analysis setup **
.DC LIN     
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "cc112.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
