* C:\Users\ASADULLAH\Documents\Schematic4.sch

* Schematics Version 9.2
* Fri Aug 18 23:31:28 2017


.PARAM         VAR=10 

** Analysis setup **
.DC LIN PARAM VAR 0 20 1 
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Schematic4.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
