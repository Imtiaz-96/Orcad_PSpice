* C:\Users\ASADULLAH\Documents\Schematic1.sch

* Schematics Version 9.2
* Sat Aug 12 23:26:48 2017



** Analysis setup **
.DC LIN V_V1 5 20 1 
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Schematic1.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
