* C:\Users\ASADULLAH\Documents\EEEex2figfour.sch

* Schematics Version 9.2
* Wed Jan 24 17:41:41 2018



** Analysis setup **
.ac DEC 20 10 100g
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "EEEex2figfour.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
