* C:\Users\ASADULLAH\Documents\chapfourfigthree.sch

* Schematics Version 9.2
* Sun Jan 28 00:38:17 2018



** Analysis setup **
.DC LIN V_Vgg 0 5 .01 
+ LIN V_Vdd 0 5 1 
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "chapfourfigthree.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
