* C:\Users\ASADULLAH\Documents\sixfourone.sch

* Schematics Version 9.2
* Mon Nov 27 11:39:16 2017



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "sixfourone.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
