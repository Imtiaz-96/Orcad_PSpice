* C:\Users\ASADULLAH\Documents\Schematic2.sch

* Schematics Version 9.2
* Tue Aug 15 23:25:32 2017



** Analysis setup **
.tran 0ns 1000ns
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Schematic2.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
