* C:\Users\ASADULLAH\Documents\sicbyone.sch

* Schematics Version 9.2
* Thu Jan 25 23:03:55 2018



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "sicbyone.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
