* C:\Users\ASADULLAH\Documents\sixaone.sch

* Schematics Version 9.2
* Sat Nov 25 12:03:11 2017



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "sixaone.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
