* C:\Users\ASADULLAH\Documents\figuresixto three.sch

* Schematics Version 9.2
* Sat Jan 27 12:25:31 2018



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "figuresixto three.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
