* C:\Users\ASADULLAH\Documents\Schematic5.sch

* Schematics Version 9.2
* Fri Aug 18 23:36:08 2017


.PARAM         VAR=10 

** Analysis setup **
.DC LIN PARAM VAR 1 20 1 
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Schematic5.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
