* C:\Users\ASADULLAH\Documents\newEEEex2figuretwo.sch

* Schematics Version 9.2
* Wed Oct 25 11:08:59 2017



** Analysis setup **
.ac DEC 20 10 100meg
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "newEEEex2figuretwo.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
