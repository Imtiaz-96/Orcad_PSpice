* C:\Users\ASADULLAH\Documents\Schematic3.sch

* Schematics Version 9.2
* Fri Aug 18 23:19:07 2017


.PARAM         RVAR=10 

** Analysis setup **
.DC LIN PARAM RVAR .1 20 .1 
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Schematic3.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
