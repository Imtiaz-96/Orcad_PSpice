* C:\Users\ASADULLAH\Documents\chapfivefigthree.sch

* Schematics Version 9.2
* Thu Jan 25 22:27:59 2018



** Analysis setup **
.ac DEC 20 10 1meg
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "chapfivefigthree.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
