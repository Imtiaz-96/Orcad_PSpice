* C:\Users\ASADULLAH\Documents\eeeextwofigurethree.sch

* Schematics Version 9.2
* Tue Jan 30 22:36:14 2018



** Analysis setup **
.ac DEC 20 10 100meg
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "eeeextwofigurethree.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
